/*
	This is our top-level module
*/
module Matrix_Multiplier(


);




endmodule 