module mux2(
	input [5:0] address,
	input reset,
	output reg [5:0] writeAddress
);

always@(*) begin
	if(reset) begin
		writeAddress = 0;
	end else begin
		writeAddress = address;
	end
end

endmodule

